module site

struct Site {

}

fn (site Site) create() ? Site {
}

fn (site Site) read() ? Site {
}

fn (site Site) update() ? Site {
}

fn (site Site) delete() ? Site {
}

pub fn create_site() {
}

pub fn read_site() {
}

pub fn update_site() {
}

pub fn delete_site() {
    function := Site.delete()
	
}