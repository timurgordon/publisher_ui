module ui_kit

import vweb
import os

pub interface Component {
	mut:
	template string
}