module ui_kit

pub struct Login {
	heading string
	login Action
	remember Action
}