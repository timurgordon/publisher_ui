module ui_kit

pub struct Login {
	pub:
	heading string
	login Action
	remember Action
}